// *********************************************************************************
// Author       : huzhengxuan
// E-mail       : huzhengxuan23s@ict.ac.cn
// File         : carry4.v
// Create       : 2023-12-05 16:55
// *********************************************************************************
// Description  : 
//                carry4
//==================================================================================
// Revision History:
// Date         By              Revision        Change Description
//----------------------------------------------------------------------------------
// 2023-12-05   huzhengxuan        1.0             Original
//==================================================================================

module carry4 
(
    input   [3:0]       p,
    input   [3:0]       g,
    input                 cin,
    output               P,G,
    output [2:0]       cout
);

assign P = &p;
assign G = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]);

assign cout[0] = g[0] | (p[0] & cin);
assign cout[1] = g[1] | (p[1] & g[0]) | (p[1] & p[0] & cin);
assign cout[2] = g[2] | (p[2] & g[1]) | (p[2] & p[1] & g[0]) | (p[2] & p[1] & p[0] & cin);

endmodule


