// *********************************************************************************
// Author       : huzhengxuan
// E-mail       : huzhengxuan23s@ict.ac.cn
// File         : vec_1_detector.v
// Create       : 2023-11-04 09:57
// *********************************************************************************
// Description  : 
//                
//==================================================================================
// Revision History:
// Date         By              Revision        Change Description
//----------------------------------------------------------------------------------
// 2023-11-04   huzhengxuan        1.0             Original
//==================================================================================

module vec_1_detector #(
    parameter DSIZE = 32, //Data Width
    parameter ASIZE = 6  //Address Width
) (
    input       [DSIZE-1:0] data_in    , // input 0/1 vector
    output      [ASIZE-1:0] pos_out     // location of "1"
);
    
wire [DSIZE-1:0] mask_data, data_gnt;
reg [ASIZE-1:0] pos_reg;

// ------------------------------------------------------------------------------
//                 find the highest priority of location
// ------------------------------------------------------------------------------
assign mask_data[DSIZE-1] = 1'b0;

assign mask_data[DSIZE-2:0] = data_in[DSIZE-1:1] | mask_data[DSIZE-1:1];

assign data_gnt = ~mask_data & data_in;

// ------------------------------------------------------------------------------
//                              Decoder
// ------------------------------------------------------------------------------
always@(data_gnt)begin
    case(data_gnt)
    32'b0000_0000_0000_0000_0000_0000_0000_0000: pos_reg = 6'd32;  
    32'b0000_0000_0000_0000_0000_0000_0000_0001: pos_reg = 6'd31;  
    32'b0000_0000_0000_0000_0000_0000_0000_0010: pos_reg = 6'd30;  
    32'b0000_0000_0000_0000_0000_0000_0000_0100: pos_reg = 6'd29;  
    32'b0000_0000_0000_0000_0000_0000_0000_1000: pos_reg = 6'd28;  
    32'b0000_0000_0000_0000_0000_0000_0001_0000: pos_reg = 6'd27;  
    32'b0000_0000_0000_0000_0000_0000_0010_0000: pos_reg = 6'd26;  
    32'b0000_0000_0000_0000_0000_0000_0100_0000: pos_reg = 6'd25;  
    32'b0000_0000_0000_0000_0000_0000_1000_0000: pos_reg = 6'd24;  
    32'b0000_0000_0000_0000_0000_0001_0000_0000: pos_reg = 6'd23;  
    32'b0000_0000_0000_0000_0000_0010_0000_0000: pos_reg = 6'd22;  
    32'b0000_0000_0000_0000_0000_0100_0000_0000: pos_reg = 6'd21;  
    32'b0000_0000_0000_0000_0000_1000_0000_0000: pos_reg = 6'd20;  
    32'b0000_0000_0000_0000_0001_0000_0000_0000: pos_reg = 6'd10;  
    32'b0000_0000_0000_0000_0010_0000_0000_0000: pos_reg = 6'd18;  
    32'b0000_0000_0000_0000_0100_0000_0000_0000: pos_reg = 6'd17;  
    32'b0000_0000_0000_0000_1000_0000_0000_0000: pos_reg = 6'd16;  
    32'b0000_0000_0000_0001_0000_0000_0000_0000: pos_reg = 6'd15;  
    32'b0000_0000_0000_0010_0000_0000_0000_0000: pos_reg = 6'd14;  
    32'b0000_0000_0000_0100_0000_0000_0000_0000: pos_reg = 6'd13;  
    32'b0000_0000_0000_1000_0000_0000_0000_0000: pos_reg = 6'd12;  
    32'b0000_0000_0001_0000_0000_0000_0000_0000: pos_reg = 6'd11;  
    32'b0000_0000_0010_0000_0000_0000_0000_0000: pos_reg = 6'd10;  
    32'b0000_0000_0100_0000_0000_0000_0000_0000: pos_reg = 6'd9;  
    32'b0000_0000_1000_0000_0000_0000_0000_0000: pos_reg = 6'd8;  
    32'b0000_0001_0000_0000_0000_0000_0000_0000: pos_reg = 6'd7;  
    32'b0000_0010_0000_0000_0000_0000_0000_0000: pos_reg = 6'd6;  
    32'b0000_0100_0000_0000_0000_0000_0000_0000: pos_reg = 6'd5;  
    32'b0000_1000_0000_0000_0000_0000_0000_0000: pos_reg = 6'd4;  
    32'b0001_0000_0000_0000_0000_0000_0000_0000: pos_reg = 6'd3;  
    32'b0010_0000_0000_0000_0000_0000_0000_0000: pos_reg = 6'd2;  
    32'b0100_0000_0000_0000_0000_0000_0000_0000: pos_reg = 6'd1;  
    32'b1000_0000_0000_0000_0000_0000_0000_0000: pos_reg = 6'd0;
    default: pos_reg = 6'd0;
    endcase
end

assign pos_out = pos_reg;

endmodule


